`include "fadd.v"

module rpfadd8(
    input cin,
    input [7:0] a,
    input [7:0] b,
    output [7:0] sum,
    output cout
);

    // TODO: write your code here

endmodule