`timescale 1ns / 1ps

module alu(
    input [7:0] a,
    input [7:0] b,
    input [2:0] opcode,
    output [7:0] result,
    output co
);

    // write your code here

endmodule