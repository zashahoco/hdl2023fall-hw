`include "bcdfadd4.v"

module bcdfadd16(
  input wire [15:0] a,
  input wire [15:0] b,
  input wire cin,
  output wire [15:0] sum,
  output wire cout
);

  // write your code here

endmodule
